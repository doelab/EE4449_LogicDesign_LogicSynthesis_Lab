library verilog;
use verilog.vl_types.all;
entity p1swtb is
end p1swtb;
