//top level file of your Lab 3