//`default_nettype none

// Starter code for Project 2.  See README.md for details

module ChipInterface
  (input  logic       CLOCK_50,
   input  logic [0:0] SW,
   input  logic [0:0] KEY,
   output logic [6:0] HEX5, HEX4, HEX3, HEX2, HEX1, HEX0);

endmodule:ChipInterface