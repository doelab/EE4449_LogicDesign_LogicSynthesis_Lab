module lfshr (clk,rst,seed,out) //16-bit linear feed back shift register
    input clk;
    input rst;
    input [15:0] seed;
    output [15:0] out;

endmodule