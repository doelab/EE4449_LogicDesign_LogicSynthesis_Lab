`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DjPctyD/U0weDUIMH5TZ9GOIik3BT/Pc9Hyeh+d26eBCUJ8Vd51TPE/jq4nOLC91
u/nT/gN60ixoTK0WqSX41dCox/Tt+yHt4bNl/djZoNfVQBFm4ji0JgUaThVdAQIX
FaijgteOUBKruoW/fO1mNNTKFEOyGWlZ1YO7e+AX46MtU90/iNrljt++1w5aB2Yc
7RFH5bUPqCc36svE1FFwAqG4kZUFcyqR1i+r0T+JDeBkGZbABCPUbbKh8hC5bmuR
g8NymRLXij6xmA2mo1CcCFH7t3iagQGaXswIdRZ/HSWf0O9AbTkoVi9VomubkyxQ
Qfxb0H410mWuPWT6/C8ZTEd61iKzDgJC636tt7QbfUE95F8NQ/onWtbmCLHhctFS
9Q2DbCNVyo8IB0PoRmt9eVr6hBlSTfM7vl/sq+Qh2qa8TFtQT5QAzx/uMYT0px0f
3z37yQX5+FwjEyxnuI98mWPYnTi4LaP1ed++FOuHIJM1wxBn3B4qBdQ4tjqOu4f1
fLuxpDisKsq4AmBItrewiOjfhVSrO1F68o0e75FZZNSNwEMKBn1XtIHu/OEf3sRT
MHkZ0JsMx77JIuYK9dIok8advbuJO2EOmjNZOWp5T2TY7V5DLWt7Dsx+xod2UfP7
aFU8tYmitltFesj5i7NM2aDcPYe2mCTktnAldEi6G3T4R4NEq3CvlNzxbVxc1c3F
hQJdU6bXUct9o19AjndmPyNDEq6dK15WXHgPuIlbNC5s4Tq+gmOYqXlkSM+4O8B5
6YqKKlfKfKOw8E4p4sd7Ijti4yi6uEqDhc8vckacBXzHZFnoJTxx0CN4f9+HPfFZ
i03IuUw4YGhf3TNSq4X6RQ5wh8dXRQW0k3PK6Ml+xqmW/WceueDtWVQW+IzLXl1q
ZjD1xTRV4dlQNx8Gx92UbdslohClvhpXrPQLZwDa60c820z/Fpex9ZxDn9/u8Kxl
fWxKwGDQ/Lv0lw7IMAVfsuQvNHAE+DOJ1heaO9A0ve0I3WyTWTxF9YdOgaHKwGM3
sQXzm+ajf0ADftchKTXA5x4xcugxkprwt5mgL0w0/hV4rQziBCxxz9rGUyhBOjZ/
8HqkQSeh1xLjayxbfpAeudv7TJBFQyAeOxuGyURr5ZcqfQIdprLrTaKMgYYtYlnZ
iw5Dn9fWW2PnOF3ggalG4Ist8S4VJdjR4tHsViUzArJPOneS1r20hyLiZU8nmt2Z
/0PT3dDJC70RQ+Ugmp8miAsmDCFLcUlKVwuDhJbgX2uik4umgRMnVwcSk1M1BJk8
agHQzSYJA7xzYbAVIXubSyROTzJP3kd8cXYcjo5UKnhyfRYKXDqrM5tO2M+Zn33S
sIe3eL7HqniOJfqlXB+zcC5HLfa3G7lXsMGVSlTewLoUj9yQJzAbuy3fVRICTKXM
iaULkgauhmc7vXgF3wAEvGooCzoUucXlCHwh3cD0hPlKQUkLMtdbxX04b9lMghsN
RWQhBFLTProLdSZyLTQrQA==
`protect END_PROTECTED
