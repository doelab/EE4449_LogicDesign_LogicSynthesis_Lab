module downstream // For Altera DE10s board
	(input	logic				clk, reset_l,
	 input	logic	done,
	 input logic [7:0] downstream_in,
     output logic [7:0] downstream_out
	 );

////////////////
//write your code here

////////////////

endmodule
