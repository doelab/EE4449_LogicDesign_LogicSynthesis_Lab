library verilog;
use verilog.vl_types.all;
entity BCDtoSevenSegmentTest is
end BCDtoSevenSegmentTest;
