module p1 // For Altera DE10s board
	(input	logic	CLOCK_50,
     input     logic     KEY0,
     input logic KEY2,
     output logic LED0,
     output logic [6:0] HEX3,HEX2, //testbench out
     output logic [6:0] HEX1,HEX0 //downstream out
     );

////////////////
//write your code here


////////////////

endmodule